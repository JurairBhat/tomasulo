/* This module gets the instruction from the memory
puts the data in instruction register */
module fetch(
  input [7:0] mem_address,
  input mem_read ,
  input ir_w , // it only write in intruction register if ir_w = 1
  output [31:0] opcode
  );

  // code to put
endmodule

module(
    input [31:0]

  )

  )
